module MIDIsampler	(
						input signal,clk,rst,
						output[7:0] LED
					);

endmodule 